module CSA_2bit (X,Y,Cin,Cout,Sum);

input 	[1:0]		X;
input 	[1:0]		Y;
input 			Cin;
output 			Cout;
output	[1:0]		Sum;



wire			S_C1;
wire			S_C0;
wire			Carry_out_C0;
wire			Carry_out_C1;
wire			Cin_select;



Full_Adder FA_LSB(
	.X(X[0]),
	.Y(Y[0]),
	.Cin(Cin),
	.Cout(Cin_select),
	.Sum(Sum[0])
);

Full_Adder FA_MSB_C0(
	.X(X[1]),
	.Y(Y[1]),
	.Cin(1'b0),
	.Cout(Carry_out_C0),
	.Sum(S_C0)
);


Full_Adder FA_MSB_C1(
	.X(X[1]),
	.Y(Y[1]),
	.Cin(1'b1),
	.Cout(Carry_out_C1),
	.Sum(S_C1)
);


assign Sum[1] = (Cin_select)? S_C1 : S_C0;
assign Cout = (Cin_select)? Carry_out_C1 : Carry_out_C0; 

endmodule	















